`timescale 1ns / 1ps

module lut(
    input clk,
	 input reset,
    input [7:0] phase,
    output [7:0] sin_out,
	 output [7:0] cos_out
    );

reg [7:0]sin_reg;
reg [7:0]cos_reg;
reg [7:0]rom[255:0];

wire [7:0]index;
wire [7:0]cos_index;

assign sin_out = sin_reg;
assign cos_out = cos_reg;

assign index = phase;
assign cos_index = phase+8'd64;

initial
begin
	//$readmemh("ram.data", rom, 0, 255);
	sin_reg = 0;
	cos_reg = 0;
	rom[0] = 8'h03;
	rom[1] = 8'h06;
	rom[2] = 8'h09;
	rom[3] = 8'h0C;
	rom[4] = 8'h10;
	rom[5] = 8'h13;
	rom[6] = 8'h16;
	rom[7] = 8'h19;
	rom[8] = 8'h1C;
	rom[9] = 8'h1F;
	rom[10] = 8'h22;
	rom[11] = 8'h25;
	rom[12] = 8'h28;
	rom[13] = 8'h2B;
	rom[14] = 8'h2E;
	rom[15] = 8'h31;
	rom[16] = 8'h33;
	rom[17] = 8'h36;
	rom[18] = 8'h39;
	rom[19] = 8'h3C;
	rom[20] = 8'h3F;
	rom[21] = 8'h41;
	rom[22] = 8'h44;
	rom[23] = 8'h47;
	rom[24] = 8'h49;
	rom[25] = 8'h4C;
	rom[26] = 8'h4E;
	rom[27] = 8'h51;
	rom[28] = 8'h53;
	rom[29] = 8'h55;
	rom[30] = 8'h58;
	rom[31] = 8'h5A;
	rom[32] = 8'h5C;
	rom[33] = 8'h5E;
	rom[34] = 8'h60;
	rom[35] = 8'h62;
	rom[36] = 8'h64;
	rom[37] = 8'h66;
	rom[38] = 8'h68;
	rom[39] = 8'h6A;
	rom[40] = 8'h6B;
	rom[41] = 8'h6D;
	rom[42] = 8'h6F;
	rom[43] = 8'h70;
	rom[44] = 8'h71;
	rom[45] = 8'h73;
	rom[46] = 8'h74;
	rom[47] = 8'h75;
	rom[48] = 8'h76;
	rom[49] = 8'h78;
	rom[50] = 8'h79;
	rom[51] = 8'h7A;
	rom[52] = 8'h7A;
	rom[53] = 8'h7B;
	rom[54] = 8'h7C;
	rom[55] = 8'h7D;
	rom[56] = 8'h7D;
	rom[57] = 8'h7E;
	rom[58] = 8'h7E;
	rom[59] = 8'h7E;
	rom[60] = 8'h7F;
	rom[61] = 8'h7F;
	rom[62] = 8'h7F;
	rom[63] = 8'h7F;
	rom[64] = 8'h7F;
	rom[65] = 8'h7F;
	rom[66] = 8'h7F;
	rom[67] = 8'h7E;
	rom[68] = 8'h7E;
	rom[69] = 8'h7E;
	rom[70] = 8'h7D;
	rom[71] = 8'h7D;
	rom[72] = 8'h7C;
	rom[73] = 8'h7B;
	rom[74] = 8'h7A;
	rom[75] = 8'h7A;
	rom[76] = 8'h79;
	rom[77] = 8'h78;
	rom[78] = 8'h76;
	rom[79] = 8'h75;
	rom[80] = 8'h74;
	rom[81] = 8'h73;
	rom[82] = 8'h71;
	rom[83] = 8'h70;
	rom[84] = 8'h6F;
	rom[85] = 8'h6D;
	rom[86] = 8'h6B;
	rom[87] = 8'h6A;
	rom[88] = 8'h68;
	rom[89] = 8'h66;
	rom[90] = 8'h64;
	rom[91] = 8'h62;
	rom[92] = 8'h60;
	rom[93] = 8'h5E;
	rom[94] = 8'h5C;
	rom[95] = 8'h5A;
	rom[96] = 8'h58;
	rom[97] = 8'h55;
	rom[98] = 8'h53;
	rom[99] = 8'h51;
	rom[100] = 8'h4E;
	rom[101] = 8'h4C;
	rom[102] = 8'h49;
	rom[103] = 8'h47;
	rom[104] = 8'h44;
	rom[105] = 8'h41;
	rom[106] = 8'h3F;
	rom[107] = 8'h3C;
	rom[108] = 8'h39;
	rom[109] = 8'h36;
	rom[110] = 8'h33;
	rom[111] = 8'h31;
	rom[112] = 8'h2E;
	rom[113] = 8'h2B;
	rom[114] = 8'h28;
	rom[115] = 8'h25;
	rom[116] = 8'h22;
	rom[117] = 8'h1F;
	rom[118] = 8'h1C;
	rom[119] = 8'h19;
	rom[120] = 8'h16;
	rom[121] = 8'h13;
	rom[122] = 8'h10;
	rom[123] = 8'h0C;
	rom[124] = 8'h09;
	rom[125] = 8'h06;
	rom[126] = 8'h03;
	rom[127] = 8'h00;
	rom[128] = 8'hFD;
	rom[129] = 8'hFA;
	rom[130] = 8'hF7;
	rom[131] = 8'hF4;
	rom[132] = 8'hF0;
	rom[133] = 8'hED;
	rom[134] = 8'hEA;
	rom[135] = 8'hE7;
	rom[136] = 8'hE4;
	rom[137] = 8'hE1;
	rom[138] = 8'hDE;
	rom[139] = 8'hDB;
	rom[140] = 8'hD8;
	rom[141] = 8'hD5;
	rom[142] = 8'hD2;
	rom[143] = 8'hCF;
	rom[144] = 8'hCD;
	rom[145] = 8'hCA;
	rom[146] = 8'hC7;
	rom[147] = 8'hC4;
	rom[148] = 8'hC1;
	rom[149] = 8'hBF;
	rom[150] = 8'hBC;
	rom[151] = 8'hB9;
	rom[152] = 8'hB7;
	rom[153] = 8'hB4;
	rom[154] = 8'hB2;
	rom[155] = 8'hAF;
	rom[156] = 8'hAD;
	rom[157] = 8'hAB;
	rom[158] = 8'hA8;
	rom[159] = 8'hA6;
	rom[160] = 8'hA4;
	rom[161] = 8'hA2;
	rom[162] = 8'hA0;
	rom[163] = 8'h9E;
	rom[164] = 8'h9C;
	rom[165] = 8'h9A;
	rom[166] = 8'h98;
	rom[167] = 8'h96;
	rom[168] = 8'h95;
	rom[169] = 8'h93;
	rom[170] = 8'h91;
	rom[171] = 8'h90;
	rom[172] = 8'h8F;
	rom[173] = 8'h8D;
	rom[174] = 8'h8C;
	rom[175] = 8'h8B;
	rom[176] = 8'h8A;
	rom[177] = 8'h88;
	rom[178] = 8'h87;
	rom[179] = 8'h86;
	rom[180] = 8'h86;
	rom[181] = 8'h85;
	rom[182] = 8'h84;
	rom[183] = 8'h83;
	rom[184] = 8'h83;
	rom[185] = 8'h82;
	rom[186] = 8'h82;
	rom[187] = 8'h82;
	rom[188] = 8'h81;
	rom[189] = 8'h81;
	rom[190] = 8'h81;
	rom[191] = 8'h81;
	rom[192] = 8'h81;
	rom[193] = 8'h81;
	rom[194] = 8'h81;
	rom[195] = 8'h82;
	rom[196] = 8'h82;
	rom[197] = 8'h82;
	rom[198] = 8'h83;
	rom[199] = 8'h83;
	rom[200] = 8'h84;
	rom[201] = 8'h85;
	rom[202] = 8'h86;
	rom[203] = 8'h86;
	rom[204] = 8'h87;
	rom[205] = 8'h88;
	rom[206] = 8'h8A;
	rom[207] = 8'h8B;
	rom[208] = 8'h8C;
	rom[209] = 8'h8D;
	rom[210] = 8'h8F;
	rom[211] = 8'h90;
	rom[212] = 8'h91;
	rom[213] = 8'h93;
	rom[214] = 8'h95;
	rom[215] = 8'h96;
	rom[216] = 8'h98;
	rom[217] = 8'h9A;
	rom[218] = 8'h9C;
	rom[219] = 8'h9E;
	rom[220] = 8'hA0;
	rom[221] = 8'hA2;
	rom[222] = 8'hA4;
	rom[223] = 8'hA6;
	rom[224] = 8'hA8;
	rom[225] = 8'hAB;
	rom[226] = 8'hAD;
	rom[227] = 8'hAF;
	rom[228] = 8'hB2;
	rom[229] = 8'hB4;
	rom[230] = 8'hB7;
	rom[231] = 8'hB9;
	rom[232] = 8'hBC;
	rom[233] = 8'hBF;
	rom[234] = 8'hC1;
	rom[235] = 8'hC4;
	rom[236] = 8'hC7;
	rom[237] = 8'hCA;
	rom[238] = 8'hCD;
	rom[239] = 8'hCF;
	rom[240] = 8'hD2;
	rom[241] = 8'hD5;
	rom[242] = 8'hD8;
	rom[243] = 8'hDB;
	rom[244] = 8'hDE;
	rom[245] = 8'hE1;
	rom[246] = 8'hE4;
	rom[247] = 8'hE7;
	rom[248] = 8'hEA;
	rom[249] = 8'hED;
	rom[250] = 8'hF0;
	rom[251] = 8'hF4;
	rom[252] = 8'hF7;
	rom[253] = 8'hFA;
	rom[254] = 8'hFD;
	rom[255] = 8'h00;
end

always @(posedge clk)
begin
	if(reset) begin
		sin_reg <= 0;
		cos_reg <= 0;
	end else begin
		sin_reg <= rom[index];
		cos_reg <= rom[cos_index];
	end
end

endmodule
